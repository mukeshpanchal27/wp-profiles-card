
<svg xmlns="http://www.w3.org/2000/svg" xmlns:xlink="http://www.w3.org/1999/xlink" version="1.1" viewBox="-10 0 532 512">
   <path fill="currentColor"
d="M256 0q70 0 128.5 34.5t93 93t34.5 128.5t-34.5 128.5t-93 93t-128.5 34.5t-128.5 -34.5t-93 -93t-34.5 -128.5t34.5 -128.5t93 -93t128.5 -34.5zM256 13q-66 0 -122 32.5t-88.5 88.5t-32.5 122t32.5 122t88.5 88.5t122 32.5t122 -32.5t88.5 -88.5t32.5 -122t-32.5 -122
t-88.5 -88.5t-122 -32.5zM256 38q59 0 109 29.5t79.5 79.5t29.5 109t-29.5 109t-79.5 79.5t-109 29.5t-109 -29.5t-79.5 -79.5t-29.5 -109t29.5 -109t79.5 -79.5t109 -29.5zM302 82q-21 0 -40 12q31 7 50.5 31.5t19.5 56.5q0 26 -14 48q26 -6 42.5 -26t16.5 -47
q0 -31 -22 -53t-53 -22zM241 108q-31 0 -53 22t-22 53t22 53t53 22t53 -22t22 -53t-22 -53t-53 -22zM350 236l-13 15q20 6 35 22q12 13 19 31q5 13 7 28l2 12h32q0 -54 -21 -82q-15 -20 -40 -25q-12 -2 -21 -1v0zM296 257l-54 53l-54 -53q-37 1 -60 22q-17 16 -25 43
q-5 20 -5 43l2 19h283q4 -36 -4 -62q-7 -23 -21 -38q-12 -12 -28 -19q-11 -5 -24 -7z" />
</svg>
